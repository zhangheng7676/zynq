module ();
    mod_name instance_name (.*);
    mod_name instance_name (.*);
endmodule